//Rudy Hill
//ECEN 2350
//Spring 2018
//
module Project2_top(CLK,KEY,SW,LED,HEX0,HEX1,HEX2,HEX3,HEX4, HEX5);
	input CLK,SW;
	input [1:0] KEY;
	output LED;
	output [7:0] HEX0,HEX1,HEX2,HEX3,HEX4,HEX5;
	wire DC_EN,DC_CLR,BCD_EN,BCD_CLR,HIGH_EN,DC_DONE,LAG;
	wire [23:0] BCD,HIGH;
	wire [10:0] Q;
	wire [7:0] DISPLAY0,DISPLAY1,DISPLAY2,DISPLAY3,DISPLAY4,DISPLAY5;
	
	Go G1(CLK,DISPLAY0,DISPLAY1,DISPLAY2,DISPLAY3,DISPLAY4,DISPLAY5);
	
	LFSR L1(LAG,Q);
	
	Down_count DO1(KEY[0],LAG,DC_EN,DC_CLR,Q,DC_DONE);
	
	High_score H1(CLK,HIGH_EN,BCD,HIGH);
	
	Clock_divider D1(CLK,LAG);
	
	FSM F1(SW,KEY,LAG,DC_DONE,DC_EN,DC_CLR,BCD_EN,BCD_CLR,HIGH_EN,LED);
	
	BCD_counter C1(BCD_EN,BCD_CLR,LAG,BCD[3:0],BCD[7:4],BCD[11:8],BCD[15:12],BCD[19:16],BCD[23:20]);
	
	BCD_decoder B1(BCD_EN,DC_CLR,CLK,SW,BCD[3:0],HIGH[3:0],HEX0,DISPLAY0);
	BCD_decoder B2(BCD_EN,DC_CLR,CLK,SW,BCD[7:4],HIGH[7:4],HEX1,DISPLAY1);
	BCD_decoder B3(BCD_EN,DC_CLR,CLK,SW,BCD[11:8],HIGH[11:8],HEX2,DISPLAY2);
	BCD_decoder B4(BCD_EN,DC_CLR,CLK,SW,BCD[15:12],HIGH[15:12],HEX3,DISPLAY3);
	BCD_decoder B5(BCD_EN,DC_CLR,CLK,SW,BCD[19:16],HIGH[19:16],HEX4,DISPLAY4);
	BCD_decoder B6(BCD_EN,DC_CLR,CLK,SW,BCD[23:20],BCD[23:20],HEX5,DISPLAY5);
endmodule

//module statemachine()

  //input button;
  //input clock;
  //input dc_done;
  //input clear;
  
  //output DC_LOAD, DC_EN, DC_CLR, BCD_EN, BCD_clear;
